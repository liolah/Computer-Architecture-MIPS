LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY pc_adder IS
  PORT (
    a : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    y : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
  );
END pc_adder;

ARCHITECTURE rtl OF pc_Adder IS
BEGIN
  PROCESS (a)
  BEGIN
    y <= a + 4;
  END PROCESS;
END rtl;
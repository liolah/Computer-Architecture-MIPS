LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY shl_2 IS
  PORT (
    x : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    y : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
  );
END shl_2;
ARCHITECTURE rtl OF shl_2 IS
BEGIN
  y(31 DOWNTO 0) <= x(29 DOWNTO 0) & "00";
END rtl;
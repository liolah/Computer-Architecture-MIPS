LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY mux_2_5bit IS
  PORT (
    a : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
    sel : IN STD_LOGIC;
    y : OUT STD_LOGIC_VECTOR(4 DOWNTO 0)
  );
END mux_2_5bit;
ARCHITECTURE rtl OF mux IS
BEGIN
  y <= a WHEN sel = '0' ELSE
    b;
END rtl;